module FA(
	input 	   x,
	input 	   y,
	input 	c_in,
	output     s, 
	output  c_out
);

/*
	Write Your Design Here ~
*/

endmodule

